module pstart_rom ( input [3:0]	addr,
						output [109:0]	data
					 );

	parameter ADDR_WIDTH = 4;
   parameter DATA_WIDTH = 110;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		  110'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 0
        110'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // 1
        110'b11111100000111111000001111111000001111100000011111000000001111111000011000110000111111110001111111000011111100, // 2 ******
        110'b01100110000011001100000110011000011000110000110001100000000110011000011100110000110110110000110011000001100110, // 3  **  **
        110'b01100110000011001100000110001000011000110000110001100000000110001000011110110000100110010000110001000001100110, // 4  **  **
        110'b01100110000011001100000110100000001100000000011000000000000110100000011111110000000110000000110100000001100110, // 5  **  **
        110'b01111100000011111000000111100000000111000000001110000000000111100000011011110000000110000000111100000001111100, // 6  *****
        110'b01100000000011011000000110100000000001100000000011000000000110100000011001110000000110000000110100000001101100, // 7  **
        110'b01100000000011001100000110000000000000110000000001100000000110000000011000110000000110000000110000000001100110, // 8  **
        110'b01100000000011001100000110001000011000110000110001100000000110001000011000110000000110000000110001000001100110, // 9  **
        110'b01100000000011001100000110011000011000110000110001100000000110011000011000110000000110000000110011000001100110, // a  **
        110'b11110000000111001100001111111000001111100000011111000000001111111000011000110000001111000001111111000011100110, // b ****
        110'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // c
        110'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // d
        110'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // e
        110'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, // f
		  };
		 
	assign data = ROM[addr];

endmodule  