module win_rom ( input [3:0]	addr,
						output [64:0]	data
					 );

	parameter ADDR_WIDTH = 4;
   parameter DATA_WIDTH = 65;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		  65'b00000000000000000000000000000000000000000000000000000000000000000, // 0
        65'b00000000000000000000000000000000000000000000000000000000000000000, // 1
        65'b11000011000011111000001100011000000110000110000011110000011000110, // 2 **    **
        65'b11000011000110001100001100011000000110000110000001100000011100110, // 3 **    **
        65'b11000011000110001100001100011000000110000110000001100000011110110, // 4 **    **
        65'b01100110000110001100001100011000000110000110000001100000011111110, // 5  **  **
        65'b00111100000110001100001100011000000110000110000001100000011011110, // 6   ****
        65'b00011000000110001100001100011000000110110110000001100000011001110, // 7    **
        65'b00011000000110001100001100011000000110110110000001100000011000110, // 8    **
        65'b00011000000110001100001100011000000111111110000001100000011000110, // 9    **
        65'b00011000000110001100001100011000000011001100000001100000011000110, // a    **
        65'b00111100000011111000000111110000000011001100000011110000011000110, // b   ****
        65'b00000000000000000000000000000000000000000000000000000000000000000, // c
        65'b00000000000000000000000000000000000000000000000000000000000000000, // d
        65'b00000000000000000000000000000000000000000000000000000000000000000, // e
        65'b00000000000000000000000000000000000000000000000000000000000000000, // f
		  };
		 
	assign data = ROM[addr];

endmodule  