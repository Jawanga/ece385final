module block_SM (input Clk,
					  input Reset,
					  