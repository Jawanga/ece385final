module title_rom ( input [3:0]	addr,
						output [40:0]	data
					 );

	parameter ADDR_WIDTH = 4;
   parameter DATA_WIDTH = 41;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
		  41'b00000000000000000000000000000000000000000, // 0
        41'b00000000000000000000000000000000000000000, // 1
        41'b11111000000110001100001111111000011111111, // 2 *****
        41'b01101100000110001100000110011000011011011, // 3  ** **
        41'b01100110000110001100000110001000010011001, // 4  **  **
        41'b01100110000110001100000110100000000011000, // 5  **  **
        41'b01100110000110001100000111100000000011000, // 6  **  **
        41'b01100110000110001100000110100000000011000, // 7  **  **
        41'b01100110000110001100000110000000000011000, // 8  **  **
        41'b01100110000110001100000110001000000011000, // 9  **  **
        41'b01101100000110001100000110011000000011000, // a  ** **
        41'b11111000000011111000001111111000000111100, // b *****
        41'b00000000000000000000000000000000000000000, // c
        41'b00000000000000000000000000000000000000000, // d
        41'b00000000000000000000000000000000000000000, // e
        41'b00000000000000000000000000000000000000000 // f
		  };
		 
	assign data = ROM[addr];

endmodule  